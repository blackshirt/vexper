module siroup






