module siroup

fn (c CPool) parse_rup(inp Rup) Rup {
	out := Rup{}
	return out
}